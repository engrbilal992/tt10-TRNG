`timescale 1ns/1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:20:19 06/03/2008 
// Design Name: 
// Module Name:    ch_xyz 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

//===========================================================================================

module ch_xyz	( 
				x,
				y,
				z,
				CH
			);

//===========================================================================================

input	[31:0]			x;
input	[31:0]			y;
input	[31:0]			z;
output	[31:0]			CH;

//===========================================================================================

assign	CH = ( (x & y) ^ ( (~x) & z) );

//--------------------------------------------------------------------------------------------------------

endmodule
